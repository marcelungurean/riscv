module Alu(
    input [31:0] io_a,
    input [31:0] io_b,
    input [3:0] io_op,
    output[31:0] io_out,
    output io_zero
);

  wire T0;
  wire T1;
  wire[31:0] alu_out;
  wire[31:0] T2;
  wire[31:0] T3;
  wire[31:0] T4;
  wire[31:0] T5;
  wire[31:0] T6;
  wire[31:0] T7;
  wire[31:0] T8;
  wire[31:0] T9;
  wire[31:0] T10;
  wire[31:0] T11;
  wire[31:0] T12;
  wire[31:0] T13;
  wire[31:0] T14;
  wire[31:0] T15;
  wire[31:0] T16;
  wire T17;
  wire[31:0] T18;
  wire[31:0] T19;
  wire[4:0] alu_shamt;
  wire[4:0] T20;
  wire[31:0] T21;
  wire T22;
  wire[31:0] T23;
  wire[31:0] T24;
  wire T25;
  wire[31:0] T26;
  wire[31:0] T27;
  wire[62:0] T28;
  wire T29;
  wire[31:0] T67;
  wire T30;
  wire T31;
  wire T32;
  wire[31:0] T68;
  wire T33;
  wire T34;
  wire[31:0] T35;
  wire[31:0] T36;
  wire T37;
  wire[31:0] T69;
  wire T38;
  wire T39;
  wire T40;
  wire[31:0] T70;
  wire T41;
  wire T42;
  wire T43;
  wire[31:0] T71;
  wire T44;
  wire T45;
  wire T46;
  wire[31:0] T72;
  wire T47;
  wire T48;
  wire[31:0] T49;
  wire[31:0] T50;
  wire T51;
  wire[31:0] T52;
  wire[31:0] T53;
  wire T54;
  wire[31:0] T55;
  wire[31:0] T56;
  wire T57;
  wire[31:0] T58;
  wire[31:0] T59;
  wire T60;
  wire[31:0] T61;
  wire[31:0] T62;
  wire T63;
  wire[31:0] T64;
  wire[31:0] T65;
  wire T66;


  assign io_zero = T0;
  assign T0 = T1 ? 1'h1 : 1'h0;
  assign T1 = io_out == 32'h0;
  assign io_out = alu_out;
  assign alu_out = T2;
  assign T2 = T66 ? T64 : T3;
  assign T3 = T63 ? T61 : T4;
  assign T4 = T60 ? T58 : T5;
  assign T5 = T57 ? T55 : T6;
  assign T6 = T54 ? T52 : T7;
  assign T7 = T51 ? T72 : T8;
  assign T8 = T46 ? T71 : T9;
  assign T9 = T43 ? T70 : T10;
  assign T10 = T40 ? T69 : T11;
  assign T11 = T37 ? T68 : T12;
  assign T12 = T32 ? T67 : T13;
  assign T13 = T29 ? T26 : T14;
  assign T14 = T25 ? T23 : T15;
  assign T15 = T22 ? T18 : T16;
  assign T16 = T17 ? io_a : 32'h0;
  assign T17 = io_op == 4'hf;
  assign T18 = T19;
  assign T19 = $signed(T21) >>> alu_shamt;
  assign alu_shamt = T20;
  assign T20 = io_b[4:0];
  assign T21 = io_a;
  assign T22 = io_op == 4'he;
  assign T23 = T24;
  assign T24 = io_a >> alu_shamt;
  assign T25 = io_op == 4'hd;
  assign T26 = T27;
  assign T27 = T28[31:0];
  assign T28 = io_a << alu_shamt;
  assign T29 = io_op == 4'hc;
  assign T67 = {31'h0, T30};
  assign T30 = T31;
  assign T31 = io_b <= io_a;
  assign T32 = io_op == 4'hb;
  assign T68 = {31'h0, T33};
  assign T33 = T34;
  assign T34 = $signed(T36) <= $signed(T35);
  assign T35 = io_a;
  assign T36 = io_b;
  assign T37 = io_op == 4'ha;
  assign T69 = {31'h0, T38};
  assign T38 = T39;
  assign T39 = io_a != io_b;
  assign T40 = io_op == 4'h9;
  assign T70 = {31'h0, T41};
  assign T41 = T42;
  assign T42 = io_a == io_b;
  assign T43 = io_op == 4'h8;
  assign T71 = {31'h0, T44};
  assign T44 = T45;
  assign T45 = io_a < io_b;
  assign T46 = io_op == 4'h7;
  assign T72 = {31'h0, T47};
  assign T47 = T48;
  assign T48 = $signed(T50) < $signed(T49);
  assign T49 = io_b;
  assign T50 = io_a;
  assign T51 = io_op == 4'h6;
  assign T52 = T53;
  assign T53 = io_a ^ io_b;
  assign T54 = io_op == 4'h5;
  assign T55 = T56;
  assign T56 = io_a | io_b;
  assign T57 = io_op == 4'h4;
  assign T58 = T59;
  assign T59 = io_a & io_b;
  assign T60 = io_op == 4'h3;
  assign T61 = T62;
  assign T62 = io_a - io_b;
  assign T63 = io_op == 4'h2;
  assign T64 = T65;
  assign T65 = io_a + io_b;
  assign T66 = io_op == 4'h1;
endmodule

