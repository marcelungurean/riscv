module Decoder(
    input [31:0] io_dec_instr,
    output io_ctl_val_inst,
    output io_ctl_rf_wen,
    output[3:0] io_ctl_br_type,
    output[1:0] io_ctl_opa_sel,
    output[1:0] io_ctl_opb_sel,
    output[3:0] io_ctl_alu_func,
    output[1:0] io_ctl_wb_sel,
    output[1:0] io_ctl_mem_func,
    output io_ctl_mem_en,
    output[2:0] io_ctl_msk_sel,
    output[2:0] io_ctl_csr_cmd
);

  wire[2:0] ctl_msk_sel;
  wire[2:0] T0;
  wire[2:0] T1;
  wire[2:0] T2;
  wire[2:0] T3;
  wire[2:0] T4;
  wire[2:0] T5;
  wire[2:0] T6;
  wire[2:0] T7;
  wire[2:0] T8;
  wire[2:0] T9;
  wire[2:0] T10;
  wire[2:0] T11;
  wire[2:0] T12;
  wire[2:0] T13;
  wire[2:0] T14;
  wire[2:0] T15;
  wire T16;
  wire[31:0] T17;
  wire T18;
  wire[31:0] T19;
  wire T20;
  wire[31:0] T21;
  wire T22;
  wire[31:0] T23;
  wire T24;
  wire[31:0] T25;
  wire T26;
  wire[31:0] T27;
  wire T28;
  wire[31:0] T29;
  wire T30;
  wire[31:0] T31;
  wire T32;
  wire[31:0] T33;
  wire T34;
  wire[31:0] T35;
  wire T36;
  wire[31:0] T37;
  wire T38;
  wire[31:0] T39;
  wire T40;
  wire[31:0] T41;
  wire T42;
  wire[31:0] T43;
  wire T44;
  wire[31:0] T45;
  wire T46;
  wire[31:0] T47;
  wire T48;
  wire[31:0] T49;
  wire ctl_mem_en;
  wire T50;
  wire T51;
  wire T52;
  wire T53;
  wire T54;
  wire T55;
  wire T56;
  wire T57;
  wire T58;
  wire T59;
  wire T60;
  wire T61;
  wire T62;
  wire T63;
  wire T64;
  wire T65;
  wire T66;
  wire[31:0] T67;
  wire[1:0] ctl_mem_func;
  wire[1:0] T68;
  wire[1:0] T69;
  wire[1:0] T70;
  wire[1:0] T71;
  wire[1:0] T72;
  wire[1:0] T73;
  wire[1:0] T74;
  wire[1:0] T75;
  wire[1:0] T76;
  wire[1:0] T77;
  wire[1:0] T78;
  wire[1:0] T79;
  wire[1:0] T80;
  wire[1:0] T81;
  wire[1:0] T82;
  wire[1:0] T83;
  wire[1:0] T84;
  wire[1:0] ctl_wb_sel;
  wire[1:0] T85;
  wire[1:0] T86;
  wire[1:0] T87;
  wire[1:0] T88;
  wire[1:0] T89;
  wire[1:0] T90;
  wire[1:0] T91;
  wire[1:0] T92;
  wire[1:0] T93;
  wire[1:0] T94;
  wire[1:0] T95;
  wire[1:0] T96;
  wire[1:0] T97;
  wire[1:0] T98;
  wire[3:0] ctl_alu_func;
  wire[3:0] T99;
  wire[3:0] T100;
  wire[3:0] T101;
  wire[3:0] T102;
  wire[3:0] T103;
  wire[3:0] T104;
  wire[3:0] T105;
  wire[3:0] T106;
  wire[3:0] T107;
  wire[3:0] T108;
  wire[3:0] T109;
  wire[3:0] T110;
  wire[3:0] T111;
  wire[3:0] T112;
  wire[3:0] T113;
  wire[3:0] T114;
  wire[3:0] T115;
  wire[3:0] T116;
  wire[3:0] T117;
  wire[3:0] T118;
  wire[3:0] T119;
  wire[3:0] T120;
  wire[3:0] T121;
  wire[3:0] T122;
  wire[3:0] T123;
  wire[3:0] T124;
  wire[3:0] T125;
  wire[3:0] T126;
  wire[3:0] T127;
  wire[3:0] T128;
  wire[3:0] T129;
  wire[3:0] T130;
  wire[3:0] T131;
  wire[3:0] T132;
  wire[3:0] T133;
  wire[3:0] T134;
  wire T135;
  wire[31:0] T136;
  wire T137;
  wire[31:0] T138;
  wire T139;
  wire[31:0] T140;
  wire T141;
  wire[31:0] T142;
  wire T143;
  wire[31:0] T144;
  wire T145;
  wire[31:0] T146;
  wire T147;
  wire[31:0] T148;
  wire T149;
  wire[31:0] T150;
  wire T151;
  wire[31:0] T152;
  wire T153;
  wire[31:0] T154;
  wire T155;
  wire[31:0] T156;
  wire T157;
  wire[31:0] T158;
  wire T159;
  wire[31:0] T160;
  wire T161;
  wire[31:0] T162;
  wire T163;
  wire[31:0] T164;
  wire T165;
  wire[31:0] T166;
  wire T167;
  wire[31:0] T168;
  wire T169;
  wire[31:0] T170;
  wire T171;
  wire[31:0] T172;
  wire[1:0] ctl_opb_sel;
  wire[1:0] T173;
  wire[1:0] T174;
  wire[1:0] T175;
  wire[1:0] T176;
  wire[1:0] T177;
  wire[1:0] T178;
  wire[1:0] T179;
  wire[1:0] T180;
  wire[1:0] T181;
  wire[1:0] T182;
  wire[1:0] T183;
  wire[1:0] T184;
  wire[1:0] T185;
  wire[1:0] T186;
  wire[1:0] T187;
  wire[1:0] T188;
  wire[1:0] T189;
  wire[1:0] T190;
  wire[1:0] T191;
  wire[1:0] T192;
  wire[1:0] T193;
  wire[1:0] T194;
  wire[1:0] T195;
  wire[1:0] T196;
  wire[1:0] T197;
  wire[1:0] T198;
  wire[1:0] T199;
  wire[1:0] T200;
  wire[1:0] T201;
  wire[1:0] T202;
  wire[1:0] T203;
  wire[1:0] T204;
  wire[1:0] T205;
  wire[1:0] T206;
  wire[1:0] T207;
  wire[1:0] T208;
  wire[1:0] ctl_opa_sel;
  wire[1:0] T209;
  wire[3:0] ctl_br_type;
  wire[3:0] T210;
  wire[3:0] T211;
  wire[3:0] T212;
  wire[3:0] T213;
  wire[3:0] T214;
  wire[3:0] T215;
  wire[3:0] T216;
  wire[3:0] T217;
  wire[3:0] T218;
  wire ctl_rf_wen;
  wire T219;
  wire T220;
  wire T221;
  wire T222;
  wire T223;
  wire T224;
  wire T225;
  wire T226;
  wire T227;
  wire T228;
  wire T229;
  wire T230;
  wire T231;
  wire T232;
  wire T233;
  wire T234;
  wire T235;
  wire T236;
  wire T237;
  wire T238;
  wire T239;
  wire T240;
  wire T241;
  wire T242;
  wire T243;
  wire T244;
  wire T245;
  wire T246;
  wire T247;
  wire T248;
  wire T249;
  wire T250;
  wire T251;
  wire T252;
  wire T253;
  wire ctl_val_inst;
  wire T254;
  wire T255;
  wire T256;
  wire T257;
  wire T258;
  wire T259;
  wire T260;
  wire T261;
  wire T262;
  wire T263;
  wire T264;
  wire T265;
  wire T266;
  wire T267;
  wire T268;
  wire T269;
  wire T270;
  wire T271;
  wire T272;
  wire T273;
  wire T274;
  wire T275;
  wire T276;
  wire T277;
  wire T278;
  wire T279;
  wire T280;
  wire T281;
  wire T282;
  wire T283;
  wire T284;
  wire T285;
  wire T286;
  wire T287;
  wire T288;


  assign io_ctl_csr_cmd = 3'h0;
  assign io_ctl_msk_sel = ctl_msk_sel;
  assign ctl_msk_sel = T48 ? 3'h2 : T0;
  assign T0 = T46 ? 3'h2 : T1;
  assign T1 = T44 ? 3'h2 : T2;
  assign T2 = T42 ? 3'h2 : T3;
  assign T3 = T40 ? 3'h2 : T4;
  assign T4 = T38 ? 3'h2 : T5;
  assign T5 = T36 ? 3'h2 : T6;
  assign T6 = T34 ? 3'h2 : T7;
  assign T7 = T32 ? 3'h2 : T8;
  assign T8 = T30 ? 3'h2 : T9;
  assign T9 = T28 ? 3'h0 : T10;
  assign T10 = T26 ? 3'h3 : T11;
  assign T11 = T24 ? 3'h1 : T12;
  assign T12 = T22 ? 3'h4 : T13;
  assign T13 = T20 ? 3'h2 : T14;
  assign T14 = T18 ? 3'h0 : T15;
  assign T15 = T16 ? 3'h1 : 3'h2;
  assign T16 = T17 == 32'h1023;
  assign T17 = io_dec_instr & 32'h707f;
  assign T18 = T19 == 32'h23;
  assign T19 = io_dec_instr & 32'h707f;
  assign T20 = T21 == 32'h2003;
  assign T21 = io_dec_instr & 32'h707f;
  assign T22 = T23 == 32'h5003;
  assign T23 = io_dec_instr & 32'h707f;
  assign T24 = T25 == 32'h1003;
  assign T25 = io_dec_instr & 32'h707f;
  assign T26 = T27 == 32'h4003;
  assign T27 = io_dec_instr & 32'h707f;
  assign T28 = T29 == 32'h3;
  assign T29 = io_dec_instr & 32'h707f;
  assign T30 = T31 == 32'h6063;
  assign T31 = io_dec_instr & 32'h707f;
  assign T32 = T33 == 32'h4063;
  assign T33 = io_dec_instr & 32'h707f;
  assign T34 = T35 == 32'h7063;
  assign T35 = io_dec_instr & 32'h707f;
  assign T36 = T37 == 32'h5063;
  assign T37 = io_dec_instr & 32'h707f;
  assign T38 = T39 == 32'h1063;
  assign T39 = io_dec_instr & 32'h707f;
  assign T40 = T41 == 32'h63;
  assign T41 = io_dec_instr & 32'h707f;
  assign T42 = T43 == 32'h67;
  assign T43 = io_dec_instr & 32'h707f;
  assign T44 = T45 == 32'h6f;
  assign T45 = io_dec_instr & 32'h7f;
  assign T46 = T47 == 32'h17;
  assign T47 = io_dec_instr & 32'h7f;
  assign T48 = T49 == 32'h37;
  assign T49 = io_dec_instr & 32'h7f;
  assign io_ctl_mem_en = ctl_mem_en;
  assign ctl_mem_en = T48 ? 1'h0 : T50;
  assign T50 = T46 ? 1'h0 : T51;
  assign T51 = T44 ? 1'h0 : T52;
  assign T52 = T42 ? 1'h0 : T53;
  assign T53 = T40 ? 1'h0 : T54;
  assign T54 = T38 ? 1'h0 : T55;
  assign T55 = T36 ? 1'h0 : T56;
  assign T56 = T34 ? 1'h0 : T57;
  assign T57 = T32 ? 1'h0 : T58;
  assign T58 = T30 ? 1'h0 : T59;
  assign T59 = T28 ? 1'h1 : T60;
  assign T60 = T26 ? 1'h1 : T61;
  assign T61 = T24 ? 1'h1 : T62;
  assign T62 = T22 ? 1'h1 : T63;
  assign T63 = T20 ? 1'h1 : T64;
  assign T64 = T18 ? 1'h1 : T65;
  assign T65 = T16 ? 1'h1 : T66;
  assign T66 = T67 == 32'h2023;
  assign T67 = io_dec_instr & 32'h707f;
  assign io_ctl_mem_func = ctl_mem_func;
  assign ctl_mem_func = T48 ? 2'h0 : T68;
  assign T68 = T46 ? 2'h0 : T69;
  assign T69 = T44 ? 2'h0 : T70;
  assign T70 = T42 ? 2'h0 : T71;
  assign T71 = T40 ? 2'h0 : T72;
  assign T72 = T38 ? 2'h0 : T73;
  assign T73 = T36 ? 2'h0 : T74;
  assign T74 = T34 ? 2'h0 : T75;
  assign T75 = T32 ? 2'h0 : T76;
  assign T76 = T30 ? 2'h0 : T77;
  assign T77 = T28 ? 2'h0 : T78;
  assign T78 = T26 ? 2'h0 : T79;
  assign T79 = T24 ? 2'h0 : T80;
  assign T80 = T22 ? 2'h0 : T81;
  assign T81 = T20 ? 2'h0 : T82;
  assign T82 = T18 ? 2'h1 : T83;
  assign T83 = T16 ? 2'h1 : T84;
  assign T84 = T66 ? 2'h1 : 2'h0;
  assign io_ctl_wb_sel = ctl_wb_sel;
  assign ctl_wb_sel = T48 ? 2'h0 : T85;
  assign T85 = T46 ? 2'h0 : T86;
  assign T86 = T44 ? 2'h2 : T87;
  assign T87 = T42 ? 2'h2 : T88;
  assign T88 = T40 ? 2'h0 : T89;
  assign T89 = T38 ? 2'h0 : T90;
  assign T90 = T36 ? 2'h0 : T91;
  assign T91 = T34 ? 2'h0 : T92;
  assign T92 = T32 ? 2'h0 : T93;
  assign T93 = T30 ? 2'h0 : T94;
  assign T94 = T28 ? 2'h3 : T95;
  assign T95 = T26 ? 2'h3 : T96;
  assign T96 = T24 ? 2'h3 : T97;
  assign T97 = T22 ? 2'h3 : T98;
  assign T98 = T20 ? 2'h3 : 2'h0;
  assign io_ctl_alu_func = ctl_alu_func;
  assign ctl_alu_func = T48 ? 4'hf : T99;
  assign T99 = T46 ? 4'h1 : T100;
  assign T100 = T44 ? 4'h0 : T101;
  assign T101 = T42 ? 4'h0 : T102;
  assign T102 = T40 ? 4'h0 : T103;
  assign T103 = T38 ? 4'h0 : T104;
  assign T104 = T36 ? 4'h0 : T105;
  assign T105 = T34 ? 4'h0 : T106;
  assign T106 = T32 ? 4'h0 : T107;
  assign T107 = T30 ? 4'h0 : T108;
  assign T108 = T28 ? 4'h1 : T109;
  assign T109 = T26 ? 4'h1 : T110;
  assign T110 = T24 ? 4'h1 : T111;
  assign T111 = T22 ? 4'h1 : T112;
  assign T112 = T20 ? 4'h1 : T113;
  assign T113 = T18 ? 4'h1 : T114;
  assign T114 = T16 ? 4'h1 : T115;
  assign T115 = T66 ? 4'h1 : T116;
  assign T116 = T171 ? 4'h1 : T117;
  assign T117 = T169 ? 4'h6 : T118;
  assign T118 = T167 ? 4'h7 : T119;
  assign T119 = T165 ? 4'h5 : T120;
  assign T120 = T163 ? 4'h4 : T121;
  assign T121 = T161 ? 4'h3 : T122;
  assign T122 = T159 ? 4'hc : T123;
  assign T123 = T157 ? 4'hd : T124;
  assign T124 = T155 ? 4'he : T125;
  assign T125 = T153 ? 4'h1 : T126;
  assign T126 = T151 ? 4'h2 : T127;
  assign T127 = T149 ? 4'hc : T128;
  assign T128 = T147 ? 4'h6 : T129;
  assign T129 = T145 ? 4'h7 : T130;
  assign T130 = T143 ? 4'h5 : T131;
  assign T131 = T141 ? 4'hd : T132;
  assign T132 = T139 ? 4'he : T133;
  assign T133 = T137 ? 4'h4 : T134;
  assign T134 = T135 ? 4'h3 : 4'h0;
  assign T135 = T136 == 32'h7033;
  assign T136 = io_dec_instr & 32'hfe00707f;
  assign T137 = T138 == 32'h6033;
  assign T138 = io_dec_instr & 32'hfe00707f;
  assign T139 = T140 == 32'h40005033;
  assign T140 = io_dec_instr & 32'hfe00707f;
  assign T141 = T142 == 32'h5033;
  assign T142 = io_dec_instr & 32'hfe00707f;
  assign T143 = T144 == 32'h4033;
  assign T144 = io_dec_instr & 32'hfe00707f;
  assign T145 = T146 == 32'h3033;
  assign T146 = io_dec_instr & 32'hfe00707f;
  assign T147 = T148 == 32'h2033;
  assign T148 = io_dec_instr & 32'hfe00707f;
  assign T149 = T150 == 32'h1033;
  assign T150 = io_dec_instr & 32'hfe00707f;
  assign T151 = T152 == 32'h40000033;
  assign T152 = io_dec_instr & 32'hfe00707f;
  assign T153 = T154 == 32'h33;
  assign T154 = io_dec_instr & 32'hfe00707f;
  assign T155 = T156 == 32'h40005013;
  assign T156 = io_dec_instr & 32'hfc00707f;
  assign T157 = T158 == 32'h5013;
  assign T158 = io_dec_instr & 32'hfc00707f;
  assign T159 = T160 == 32'h1013;
  assign T160 = io_dec_instr & 32'hfc00707f;
  assign T161 = T162 == 32'h7013;
  assign T162 = io_dec_instr & 32'h707f;
  assign T163 = T164 == 32'h6013;
  assign T164 = io_dec_instr & 32'h707f;
  assign T165 = T166 == 32'h4013;
  assign T166 = io_dec_instr & 32'h707f;
  assign T167 = T168 == 32'h3013;
  assign T168 = io_dec_instr & 32'h707f;
  assign T169 = T170 == 32'h2013;
  assign T170 = io_dec_instr & 32'h707f;
  assign T171 = T172 == 32'h13;
  assign T172 = io_dec_instr & 32'h707f;
  assign io_ctl_opb_sel = ctl_opb_sel;
  assign ctl_opb_sel = T48 ? 2'h0 : T173;
  assign T173 = T46 ? 2'h1 : T174;
  assign T174 = T44 ? 2'h0 : T175;
  assign T175 = T42 ? 2'h2 : T176;
  assign T176 = T40 ? 2'h0 : T177;
  assign T177 = T38 ? 2'h0 : T178;
  assign T178 = T36 ? 2'h0 : T179;
  assign T179 = T34 ? 2'h0 : T180;
  assign T180 = T32 ? 2'h0 : T181;
  assign T181 = T30 ? 2'h0 : T182;
  assign T182 = T28 ? 2'h2 : T183;
  assign T183 = T26 ? 2'h2 : T184;
  assign T184 = T24 ? 2'h2 : T185;
  assign T185 = T22 ? 2'h2 : T186;
  assign T186 = T20 ? 2'h2 : T187;
  assign T187 = T18 ? 2'h3 : T188;
  assign T188 = T16 ? 2'h3 : T189;
  assign T189 = T66 ? 2'h3 : T190;
  assign T190 = T171 ? 2'h2 : T191;
  assign T191 = T169 ? 2'h2 : T192;
  assign T192 = T167 ? 2'h2 : T193;
  assign T193 = T165 ? 2'h2 : T194;
  assign T194 = T163 ? 2'h2 : T195;
  assign T195 = T161 ? 2'h2 : T196;
  assign T196 = T159 ? 2'h2 : T197;
  assign T197 = T157 ? 2'h2 : T198;
  assign T198 = T155 ? 2'h2 : T199;
  assign T199 = T153 ? 2'h2 : T200;
  assign T200 = T151 ? 2'h2 : T201;
  assign T201 = T149 ? 2'h2 : T202;
  assign T202 = T147 ? 2'h2 : T203;
  assign T203 = T145 ? 2'h2 : T204;
  assign T204 = T143 ? 2'h2 : T205;
  assign T205 = T141 ? 2'h2 : T206;
  assign T206 = T139 ? 2'h2 : T207;
  assign T207 = T137 ? 2'h2 : T208;
  assign T208 = T135 ? 2'h2 : 2'h0;
  assign io_ctl_opa_sel = ctl_opa_sel;
  assign ctl_opa_sel = T48 ? 2'h1 : T209;
  assign T209 = T46 ? 2'h1 : 2'h0;
  assign io_ctl_br_type = ctl_br_type;
  assign ctl_br_type = T48 ? 4'h0 : T210;
  assign T210 = T46 ? 4'h0 : T211;
  assign T211 = T44 ? 4'h7 : T212;
  assign T212 = T42 ? 4'h8 : T213;
  assign T213 = T40 ? 4'h1 : T214;
  assign T214 = T38 ? 4'h2 : T215;
  assign T215 = T36 ? 4'h3 : T216;
  assign T216 = T34 ? 4'h4 : T217;
  assign T217 = T32 ? 4'h5 : T218;
  assign T218 = T30 ? 4'h6 : 4'h0;
  assign io_ctl_rf_wen = ctl_rf_wen;
  assign ctl_rf_wen = T48 ? 1'h1 : T219;
  assign T219 = T46 ? 1'h1 : T220;
  assign T220 = T44 ? 1'h1 : T221;
  assign T221 = T42 ? 1'h1 : T222;
  assign T222 = T40 ? 1'h0 : T223;
  assign T223 = T38 ? 1'h0 : T224;
  assign T224 = T36 ? 1'h0 : T225;
  assign T225 = T34 ? 1'h0 : T226;
  assign T226 = T32 ? 1'h0 : T227;
  assign T227 = T30 ? 1'h0 : T228;
  assign T228 = T28 ? 1'h1 : T229;
  assign T229 = T26 ? 1'h1 : T230;
  assign T230 = T24 ? 1'h1 : T231;
  assign T231 = T22 ? 1'h1 : T232;
  assign T232 = T20 ? 1'h1 : T233;
  assign T233 = T18 ? 1'h0 : T234;
  assign T234 = T16 ? 1'h0 : T235;
  assign T235 = T66 ? 1'h0 : T236;
  assign T236 = T171 ? 1'h1 : T237;
  assign T237 = T169 ? 1'h1 : T238;
  assign T238 = T167 ? 1'h1 : T239;
  assign T239 = T165 ? 1'h1 : T240;
  assign T240 = T163 ? 1'h1 : T241;
  assign T241 = T161 ? 1'h1 : T242;
  assign T242 = T159 ? 1'h1 : T243;
  assign T243 = T157 ? 1'h1 : T244;
  assign T244 = T155 ? 1'h1 : T245;
  assign T245 = T153 ? 1'h1 : T246;
  assign T246 = T151 ? 1'h1 : T247;
  assign T247 = T149 ? 1'h1 : T248;
  assign T248 = T147 ? 1'h1 : T249;
  assign T249 = T145 ? 1'h1 : T250;
  assign T250 = T143 ? 1'h1 : T251;
  assign T251 = T141 ? 1'h1 : T252;
  assign T252 = T139 ? 1'h1 : T253;
  assign T253 = T137 ? 1'h1 : T135;
  assign io_ctl_val_inst = ctl_val_inst;
  assign ctl_val_inst = T48 ? 1'h1 : T254;
  assign T254 = T46 ? 1'h1 : T255;
  assign T255 = T44 ? 1'h1 : T256;
  assign T256 = T42 ? 1'h1 : T257;
  assign T257 = T40 ? 1'h1 : T258;
  assign T258 = T38 ? 1'h1 : T259;
  assign T259 = T36 ? 1'h1 : T260;
  assign T260 = T34 ? 1'h1 : T261;
  assign T261 = T32 ? 1'h1 : T262;
  assign T262 = T30 ? 1'h1 : T263;
  assign T263 = T28 ? 1'h1 : T264;
  assign T264 = T26 ? 1'h1 : T265;
  assign T265 = T24 ? 1'h1 : T266;
  assign T266 = T22 ? 1'h1 : T267;
  assign T267 = T20 ? 1'h1 : T268;
  assign T268 = T18 ? 1'h1 : T269;
  assign T269 = T16 ? 1'h1 : T270;
  assign T270 = T66 ? 1'h1 : T271;
  assign T271 = T171 ? 1'h1 : T272;
  assign T272 = T169 ? 1'h1 : T273;
  assign T273 = T167 ? 1'h1 : T274;
  assign T274 = T165 ? 1'h1 : T275;
  assign T275 = T163 ? 1'h1 : T276;
  assign T276 = T161 ? 1'h1 : T277;
  assign T277 = T159 ? 1'h1 : T278;
  assign T278 = T157 ? 1'h1 : T279;
  assign T279 = T155 ? 1'h1 : T280;
  assign T280 = T153 ? 1'h1 : T281;
  assign T281 = T151 ? 1'h1 : T282;
  assign T282 = T149 ? 1'h1 : T283;
  assign T283 = T147 ? 1'h1 : T284;
  assign T284 = T145 ? 1'h1 : T285;
  assign T285 = T143 ? 1'h1 : T286;
  assign T286 = T141 ? 1'h1 : T287;
  assign T287 = T139 ? 1'h1 : T288;
  assign T288 = T137 ? 1'h1 : T135;
endmodule

